<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 21.0.0, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<svg version="1.1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
	 viewBox="0 0 100 100" style="enable-background:new 0 0 100 100;" xml:space="preserve">
<style type="text/css">
	.st0{fill:none;stroke:#C0BFBF;stroke-width:6;stroke-miterlimit:10;}
	.st1{fill:none;stroke:#C0BFBF;stroke-width:4;stroke-miterlimit:10;}
	.st2{fill:#C0BFBF;}
	.st3{fill:none;stroke:#C0BFBF;stroke-width:6.4888;stroke-miterlimit:10;}
	.st4{fill:none;stroke:#C0BFBF;stroke-width:6.3232;stroke-miterlimit:10;}
	.st5{fill:none;stroke:#C0BFBF;stroke-width:6.3178;stroke-miterlimit:10;}
	.st6{fill:none;stroke:#C0BFBF;stroke-width:6.2472;stroke-miterlimit:10;}
	.st7{fill:none;stroke:#C0BFBF;stroke-width:6.3124;stroke-miterlimit:10;}
	.st8{fill:none;stroke:#C0BFBF;stroke-width:5;stroke-miterlimit:10;}
	.st9{fill:none;stroke:#C0BFBF;stroke-width:6.2572;stroke-miterlimit:10;}
	.st10{fill:none;stroke:#C0BFBF;stroke-width:7.4898;stroke-miterlimit:10;}
	.st11{fill:none;stroke:#C0BFBF;stroke-width:6.8128;stroke-miterlimit:10;}
	.st12{fill:none;stroke:#C0BFBF;stroke-width:6.958;stroke-miterlimit:10;}
	.st13{fill:none;stroke:#C0BFBF;stroke-width:6.9644;stroke-miterlimit:10;}
	.st14{fill:none;stroke:#C0BFBF;stroke-width:6.976;stroke-miterlimit:10;}
	.st15{fill:none;stroke:#ED2224;stroke-width:6;stroke-miterlimit:10;}
	.st16{fill:none;stroke:#ED2224;stroke-width:4;stroke-miterlimit:10;}
	.st17{fill:none;stroke:#000000;stroke-width:6;stroke-miterlimit:10;}
	.st18{fill:none;stroke:#000000;stroke-width:4;stroke-miterlimit:10;}
	.st19{font-family:'Arial-BoldMT';}
	.st20{font-size:12px;}
</style>
<g id="shadow">
	<g id="XMLID_25_">
		<g>
			<polyline class="st1" points="53.1,52.4 59,41.1 64.8,52.4 71.9,35.4 			"/>
			<g>
				<polygon class="st2" points="75.1,38 74.1,30.1 67.7,34.9 				"/>
			</g>
		</g>
	</g>
	<g id="XMLID_23_">
		<g>
			<polyline class="st1" points="47,52.4 41.1,41.1 35.3,52.4 28.2,35.4 			"/>
			<g>
				<polygon class="st2" points="32.4,34.9 26,30.1 25,38 				"/>
			</g>
		</g>
	</g>
	<line id="XMLID_329_" class="st0" x1="53" y1="5" x2="53" y2="50.5"/>
	<polygon id="XMLID_328_" class="st0" points="50,50.5 20.7,92 79.4,92 	"/>
	<line id="XMLID_327_" class="st0" x1="40.1" y1="19" x2="60.1" y2="19"/>
</g>
<g id="main">
	<g id="XMLID_21_">
		<g>
			<polyline class="st18" points="53.1,48.2 58.7,36.6 64.6,47.7 70.1,34.3 			"/>
			<g>
				<polygon points="73.4,36.9 72.3,29 66,33.8 				"/>
			</g>
		</g>
	</g>
	<g id="XMLID_16_">
		<g>
			<polyline class="st18" points="47,48.2 41.4,36.6 35.6,47.7 30,34.3 			"/>
			<g>
				<polygon points="34.1,33.8 27.8,29 26.8,36.9 				"/>
			</g>
		</g>
	</g>
	<polygon id="XMLID_325_" class="st17" points="50,45 15,95 85,95 	"/>
	<line id="XMLID_324_" class="st17" x1="50" y1="5" x2="50" y2="45"/>
	<line id="XMLID_323_" class="st18" x1="40" y1="17.2" x2="60" y2="17.2"/>
</g>
</svg>
